`timescale 1ns / 1ps

`include "xdefs.vh"

module xaddr_extdecoder_tb;