`timescale 1ns / 1ps

`include "xdefs.vh"

module xdisplay_tb;